`define CLOCK_UP `ON

`define ON  1
`define OFF 0